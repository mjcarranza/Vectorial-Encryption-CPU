module sumador(
	input [11:0] A,
	input [11:0] B,
	output [11:0] C
	);
	
	
	assign C = A + B;
	
endmodule